#top level here
